module Design3(output out, input in);

endmodule
# ECE3740_Design3
